module Adder(
  input  [31:0] io_in1,
  output [31:0] io_out
);
  assign io_out = 32'h1 + io_in1; // @[Adder.scala 13:22]
endmodule
module Register(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_; // @[Register.scala 11:23]
  assign io_out = reg_; // @[Register.scala 13:12]
  always @(posedge clock) begin
    if (reset) begin // @[Register.scala 11:23]
      reg_ <= 32'h0; // @[Register.scala 11:23]
    end else begin
      reg_ <= io_in; // @[Register.scala 12:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_ = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Count100(
  input         clock,
  input         reset,
  output [31:0] io_out
);
  wire [31:0] adder_io_in1; // @[Count100.scala 10:23]
  wire [31:0] adder_io_out; // @[Count100.scala 10:23]
  wire  register_clock; // @[Count100.scala 11:26]
  wire  register_reset; // @[Count100.scala 11:26]
  wire [31:0] register_io_in; // @[Count100.scala 11:26]
  wire [31:0] register_io_out; // @[Count100.scala 11:26]
  Adder adder ( // @[Count100.scala 10:23]
    .io_in1(adder_io_in1),
    .io_out(adder_io_out)
  );
  Register register ( // @[Count100.scala 11:26]
    .clock(register_clock),
    .reset(register_reset),
    .io_in(register_io_in),
    .io_out(register_io_out)
  );
  assign io_out = register_io_out; // @[Count100.scala 20:12]
  assign adder_io_in1 = register_io_out; // @[Count100.scala 15:18]
  assign register_clock = clock;
  assign register_reset = reset;
  assign register_io_in = register_io_out == 32'h63 ? 32'h0 : adder_io_out; // @[Count100.scala 18:19]
endmodule
